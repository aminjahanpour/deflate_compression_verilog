
            

endmodule


            